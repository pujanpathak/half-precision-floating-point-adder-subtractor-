parameter [7:0] CHAR_BLANK = 8'b00100000;

parameter [7:0] CHAR_EXCLAMATION = 8'b00100001;

parameter [7:0] CHAR_QUOTATION = 8'b00100010;

parameter [7:0] CHAR_NUMBER = 8'b00100011;

parameter [7:0] CHAR_DOLLAR = 8'b00100100;

parameter [7:0] CHAR_PERCENT = 8'b00100101;

parameter [7:0] CHAR_AMPERSAND = 8'b00100110;

parameter [7:0] CHAR_APOSTROPHE = 8'b00100111;

parameter [7:0] CHAR_LEFT_PARENTHESIS = 8'b00101000;

parameter [7:0] CHAR_RIGHT_PARENTHESIS = 8'b00101001;

parameter [7:0] CHAR_ASTERISK = 8'b00101010;

parameter [7:0] CHAR_PLUS = 8'b00101011;

parameter [7:0] CHAR_COMMA = 8'b00101100;

parameter [7:0] CHAR_HYPHEN_MINUS = 8'b00101101;

parameter [7:0] CHAR_PERIOD = 8'b00101110;

parameter [7:0] CHAR_SLASH = 8'b00101111;

parameter [7:0] CHAR_0 = 8'b00110000;

parameter [7:0] CHAR_1 = 8'b00110001;

parameter [7:0] CHAR_2 = 8'b00110010;

parameter [7:0] CHAR_3 = 8'b00110011;

parameter [7:0] CHAR_4 = 8'b00110100;

parameter [7:0] CHAR_5 = 8'b00110101;

parameter [7:0] CHAR_6 = 8'b00110110;

parameter [7:0] CHAR_7 = 8'b00110111;

parameter [7:0] CHAR_8 = 8'b00111000;

parameter [7:0] CHAR_9 = 8'b00111001;

parameter [7:0] CHAR_COLON = 8'b00111010;

parameter [7:0] CHAR_SEMICOLON = 8'b00111011;

parameter [7:0] CHAR_LESSTHAN = 8'b00111100;

parameter [7:0] CHAR_EQUALS = 8'b00111101;

parameter [7:0] CHAR_GREATERTHAN = 8'b00111110;

parameter [7:0] CHAR_QUESTION = 8'b00111111;

parameter [7:0] CHAR_AT = 8'b01000000;

parameter [7:0] CHAR_CAPITAL_A = 8'b01000001;

parameter [7:0] CHAR_CAPITAL_B = 8'b01000010;

parameter [7:0] CHAR_CAPITAL_C = 8'b01000011;

parameter [7:0] CHAR_CAPITAL_D = 8'b01000100;

parameter [7:0] CHAR_CAPITAL_E = 8'b01000101;

parameter [7:0] CHAR_CAPITAL_F = 8'b01000110;

parameter [7:0] CHAR_CAPITAL_G = 8'b01000111;

parameter [7:0] CHAR_CAPITAL_H = 8'b01001000;

parameter [7:0] CHAR_CAPITAL_I = 8'b01001001;

parameter [7:0] CHAR_CAPITAL_J = 8'b01001010;

parameter [7:0] CHAR_CAPITAL_K = 8'b01001011;

parameter [7:0] CHAR_CAPITAL_L = 8'b01001100;

parameter [7:0] CHAR_CAPITAL_M = 8'b01001101;

parameter [7:0] CHAR_CAPITAL_N = 8'b01001110;

parameter [7:0] CHAR_CAPITAL_O = 8'b01001111;

parameter [7:0] CHAR_CAPITAL_P = 8'b01010000;

parameter [7:0] CHAR_CAPITAL_Q = 8'b01010001;

parameter [7:0] CHAR_CAPITAL_R = 8'b01010010;

parameter [7:0] CHAR_CAPITAL_S = 8'b01010011;

parameter [7:0] CHAR_CAPITAL_T = 8'b01010100;

parameter [7:0] CHAR_CAPITAL_U = 8'b01010101;

parameter [7:0] CHAR_CAPITAL_V = 8'b01010110;

parameter [7:0] CHAR_CAPITAL_W = 8'b01010111;

parameter [7:0] CHAR_CAPITAL_X = 8'b01011000;

parameter [7:0] CHAR_CAPITAL_Y = 8'b01011001;

parameter [7:0] CHAR_CAPITAL_Z = 8'b01011010;

parameter [7:0] CHAR_LEFT_SQUARE_BRACKET = 8'b01011011;

parameter [7:0] CHAR_YEN = 8'b01011100;

parameter [7:0] CHAR_RIGHT_SQUARE_BRACKET = 8'b01011101;

parameter [7:0] CHAR_CIRCUMFLEX = 8'b01011110;

parameter [7:0] CHAR_LOW_LINE = 8'b01011111;

parameter [7:0] CHAR_GRAVE = 8'b01100000;

parameter [7:0] CHAR_SMALL_A = 8'b01100001;

parameter [7:0] CHAR_SMALL_B = 8'b01100010;

parameter [7:0] CHAR_SMALL_C = 8'b01100011;

parameter [7:0] CHAR_SMALL_D = 8'b01100100;

parameter [7:0] CHAR_SMALL_E = 8'b01100101;

parameter [7:0] CHAR_SMALL_F = 8'b01100110;

parameter [7:0] CHAR_SMALL_G = 8'b01100111;

parameter [7:0] CHAR_SMALL_H = 8'b01101000;

parameter [7:0] CHAR_SMALL_I = 8'b01101001;

parameter [7:0] CHAR_SMALL_J = 8'b01101010;

parameter [7:0] CHAR_SMALL_K = 8'b01101011;

parameter [7:0] CHAR_SMALL_L = 8'b01101100;

parameter [7:0] CHAR_SMALL_M = 8'b01101101;

parameter [7:0] CHAR_SMALL_N = 8'b01101110;

parameter [7:0] CHAR_SMALL_0 = 8'b01101111;

parameter [7:0] CHAR_SMALL_P = 8'b01110000;

parameter [7:0] CHAR_SMALL_Q = 8'b01110001;

parameter [7:0] CHAR_SMALL_R = 8'b01110010;

parameter [7:0] CHAR_SMALL_S = 8'b01110011;

parameter [7:0] CHAR_SMALL_T = 8'b01110100;

parameter [7:0] CHAR_SMALL_U = 8'b01110101;

parameter [7:0] CHAR_SMALL_V = 8'b01110110;

parameter [7:0] CHAR_SMALL_W = 8'b01110111;

parameter [7:0] CHAR_SMALL_X = 8'b01111000;

parameter [7:0] CHAR_SMALL_Y = 8'b01111001;

parameter [7:0] CHAR_SMALL_Z = 8'b01111010;

parameter [7:0] CHAR_LEFT_CURLY_BRACKET = 8'b01111011;

parameter [7:0] CHAR_VERTICAL_BAR = 8'b01111100;

parameter [7:0] CHAR_RIGHT_CURLY_BRACKET = 8'b01111101;

parameter [7:0] CHAR_RIGHT_ARROW = 8'b01111110;

parameter [7:0] CHAR_LEFT_ARROW = 8'b01111111;

parameter [7:0] CHAR_DIVISION = 8'b11111101;

parameter [7:0] CHAR_BLOCK = 8'b11111111;
